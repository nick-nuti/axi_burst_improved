
// SIGNALS NOT CURRENTLY USED:
    // AXI-ID   : ARID->RID, AWID->BID , identifies transaction so responses can be matched to the requester. This is for if a master allows queuing of multiple outstanding bursts
    // LOCK     : AWLOCK/ARLOCK , locked transactions (exclusive)
    // QOS      : AWQOS/ARQOS , priority hint for arbiter
    // REGION   : AWREGION/ARREGION , extra routing bits for complex interconnects
    // CACHE + PROT , cacheability and protection hints, usually for DMA/master

// FUTURE REQUIREMENTS
    // command fifo: {awid, awaddr, awlen, awsize, awburst, awprot, awcache, awqos, awregion}
    // data fifo: {wdata, wstrb}
    // resp fifo: {bresp, bid}

    // misaligned addr adjustment
    // narrow burst: yes, if someone changes AWSIZE at somepoint then keep the data_w size the same and just use write strobe accordingly
        // only allow this for AXI3

    // maybe use ID, lock, QoS, cache, prot

    // BURST type: wrapping, fixed
    
    // AWUSER, WUSER, BUSER, ARUSER, RUSER

    // with ID support "number outstanding R/W"

module axi_burst_master #(
// IP enables
    parameter WRITE_EN          =1,
    parameter READ_EN           =1,
// AXI definitions
    parameter ADDR_W            =32,
    parameter DATA_W            =64,
    // AXI
    parameter LEN_W             = 8,
    parameter LOCK_W            = 1,
    parameter QOS_W             = 4,
    parameter CACHE_W           = 4,
    parameter ABURST_W          = 2,
    parameter PROT_W            = 3,
    parameter RESP_W            = 2,
    parameter REGION_W          = 4,
    parameter ID_W              = 0,

// IP specific definitions
    parameter PAGE_SIZE_BYTES       = 4096,
    parameter SPLIT_PAGE_BOUNDARY   = 0, // 0: end burst at page boundary, >0: split burst at page boundary
    parameter BURST_POLICY          = 0, // 0: (safe) require full burst upfront, 1: stream, wait until data is present by lowering wvalid, 2: pad with dummy data if fifo empty
    parameter MISALIGN_ADJUST       = 0, // 0: disallow (results in error), >0: allow
    parameter ID_CHECK              = 0  // 0: id checking error disabled, >0: id checking error enabled
)
(
    m_axi_awaddr,
    m_axi_awprot,
    m_axi_awvalid,
    m_axi_awready,
    m_axi_awsize,
    m_axi_awburst,
    m_axi_awcache,
    m_axi_awlen,
    m_axi_awlock,
    m_axi_awqos,
    m_axi_awregion,
    m_axi_awid,
    m_axi_wdata,
    m_axi_wstrb,
    m_axi_wvalid,
    m_axi_wready,
    m_axi_wlast,
    m_axi_bresp,
    m_axi_bvalid,
    m_axi_bready,
    m_axi_bid,
    m_axi_araddr,
    m_axi_arprot,
    m_axi_arvalid,
    m_axi_arready,
    m_axi_arsize,
    m_axi_arburst,
    m_axi_arcache,
    m_axi_arlen,
    m_axi_arlock,
    m_axi_arqos,
    m_axi_arregion,
    m_axi_arid,
    m_axi_rready,
    m_axi_rdata,
    m_axi_rvalid,
    m_axi_rlast,
    m_axi_rid,
    m_axi_rresp,

    aclk,
    aresetn,

    user_w_start,
    user_w_free,

    user_w_addr,
    user_w_len,
    user_w_awsize,
    user_w_awid,

    user_w_strb,
    user_w_data,

    user_w_wready,
    user_w_wvalid,

    user_w_bid,
    user_w_status,

    user_w_bvalid,
    user_w_bready,

    user_w_cmd_error,
    user_w_underrun_event,

    user_w_data_fifo_cnt,
    user_w_data_fifo_empty,
    //user_w_data_pop_req,

    user_r_start,
    user_r_len,
    user_r_addr,
    user_r_status,
    user_r_free,
    user_r_data,
    user_r_fifo_cnt,
    user_r_fifo_full,
    user_r_data_push_req
);
    // General
    localparam BYTE = 8;
    localparam PAGE_SIZE_BYTES_CLOG = $clog2(PAGE_SIZE_BYTES);
    localparam DATA_W_CLOG = $clog2(DATA_W);
    localparam DATA_W_BYTES = DATA_W/BYTE;
    localparam DATA_W_BYTES_CLOG = $clog2(DATA_W_BYTES);
    localparam STRB_W_CLOG = $clog2(DATA_W_BYTES);

    // AXI
    localparam STRB_W           = DATA_W_BYTES;
    localparam ASIZE_W          = DATA_W_BYTES_CLOG;
    localparam MAX_BURST_BEATS  = 1 << (LEN_W);

// PORT DECLARATION
/**************** Write Address Channel Signals ****************/
    output reg [ADDR_W-1:0]             m_axi_awaddr;    // address
    output reg [PROT_W-1:0]             m_axi_awprot;    // protection - privilege and securit level of transaction
    output reg                          m_axi_awvalid;   //
    input  logic                         m_axi_awready;   //
    output reg [ASIZE_W-1:0]            m_axi_awsize;    //3'b100, // burst size - size of each transfer in the burst 3'b100 for 16 bytes/ 128 bit
    output reg [ABURST_W-1:0]           m_axi_awburst;   // fixed burst = 00, incremental = 01, wrapped burst = 10
    output reg [CACHE_W-1:0]            m_axi_awcache;   // cache type - how transaction interacts with caches
    output reg [LEN_W-1:0]              m_axi_awlen;    // number of data transfers in the burst (0-255) (done)
    output reg [LOCK_W-1:0]             m_axi_awlock;    // lock type - indicates if transaction is part of locked sequence
    output reg [QOS_W-1:0]              m_axi_awqos;     // quality of service - transaction indication of priority level
    output reg [REGION_W-1:0]           m_axi_awregion;  // region identifier - identifies targetted region
    output reg [ID_W-1:0]               m_axi_awid;
/**************** Write Data Channel Signals ****************/
    output reg [DATA_W-1:0]             m_axi_wdata;     //
    output reg [STRB_W-1:0]             m_axi_wstrb;     //
    output reg                          m_axi_wvalid;    // set to 1 when data is ready to be transferred (done)
    input  logic                         m_axi_wready;    // 
    output reg                          m_axi_wlast;     // if awlen=0 then set wlast (done)
/**************** Write Response Channel Signals ****************/
    input  logic [RESP_W-1:0]            m_axi_bresp;     // write response - status of the write transaction (00 = okay, 01 = exokay, 10 = slverr, 11 = decerr)
    input  logic                         m_axi_bvalid;    // write response valid - 0 = response not valid, 1 = response is valid
    output reg                           m_axi_bready;    // write response ready - 0 = not ready, 1 = ready
    input  logic [ID_W-1:0]              m_axi_bid;
/**************** Read Address Channel Signals ****************/
    output reg [ADDR_W-1:0]             m_axi_araddr;    // read address
    output reg [PROT_W-1:0]             m_axi_arprot;    // protection - privilege and securit level of transaction
    output reg                          m_axi_arvalid;   // 
    input  logic                        m_axi_arready;   // 
    output reg [ASIZE_W-1:0]            m_axi_arsize;    //3'b100, // burst beat size - size of each transfer in the burst 3'b100 for 16 bytes/ 128 bit
    output reg [ABURST_W-1:0]           m_axi_arburst;   // fixed burst = 00, incremental = 01, wrapped burst = 10
    output reg [CACHE_W-1:0]            m_axi_arcache;   // cache type - how transaction interacts with caches
    output reg [LEN_W-1:0]              m_axi_arlen;     // number of data transfers in the burst (0-255) (done)
    output reg [LOCK_W-1:0]             m_axi_arlock;    // lock type - indicates if transaction is part of locked sequence
    output reg [QOS_W-1:0]              m_axi_arqos;     // quality of service - transaction indication of priority level
    output reg [REGION_W-1:0]           m_axi_arregion;  // region identifier - identifies targetted region
    output reg [ID_W-1:0]               m_axi_arid;
/**************** Read Data Channel Signals ****************/
    output reg                          m_axi_rready;    // read ready - 0 = not ready, 1 = ready
    input  logic [DATA_W-1:0]            m_axi_rdata;     // 
    input  logic                         m_axi_rvalid;    // read response valid - 0 = response not valid, 1 = response is valid
    input  logic                         m_axi_rlast;     // =1 when on last read
    input  logic [ID_W-1:0]              m_axi_rid;
/**************** Read Response Channel Signals ****************/
    input  logic [RESP_W-1:0]            m_axi_rresp;     // read response - status of the read transaction (00 = okay, 01 = exokay, 10 = slverr, 11 = decerr)
/**************** System Signals ****************/
    input logic                          aclk;
    input logic                          aresetn; 
/**************** User Control Signals ****************/
//write cmd
    input  logic                         user_w_start;
    output logic                         user_w_free;
//write address
    input  logic [ADDR_W-1:0]            user_w_addr;
    input  logic [LEN_W-1:0]             user_w_len;
    input  logic [ASIZE_W-1:0]           user_w_awsize;
    input  logic [ID_W-1:0]              user_w_awid;
//write data
    input  logic [STRB_W-1:0]            user_w_strb;
    input  logic [DATA_W-1:0]            user_w_data;
//write data FIFO req/ack
    output logic                         user_w_wready; // req
    input  logic                         user_w_wvalid; // ack
//write response
    output logic [ID_W-1:0]              user_w_bid;
    output logic [RESP_W-1:0]            user_w_status; // 00:OKAY, 01:EXOKAY, 10:SLVERR, 11:DECERR
//write data req/ack
    output logic                         user_w_bvalid; // req
    input  logic                         user_w_bready; // ack
//write error
    output logic [3:0]                   user_w_cmd_error; // 00:OKAY, 01:NOROOM (1 beat can't fit before next page boundary), 
    output logic                         user_w_underrun_event;
//write fifo
    input  logic [LEN_W:0]               user_w_data_fifo_cnt; // increased the size by 1...
    input  logic                         user_w_data_fifo_empty;
    //output logic                         user_w_data_pop_req;
//read cmd
    input  logic                         user_r_start;
    input  logic [LEN_W-1:0]             user_r_len;
    input  logic [ADDR_W-1:0]            user_r_addr;
    output logic [RESP_W-1:0]            user_r_status;
    output logic                         user_r_free;
//read response
    output logic [DATA_W-1:0]            user_r_data;
//read fifo
    input  logic [LEN_W-1:0]             user_r_fifo_cnt;
    input  logic                         user_r_fifo_full;
    output reg                           user_r_data_push_req;
/*******************************************************/

// AXI W ---------------------------------------------------
generate
    if(WRITE_EN)
    begin

        logic                   start_write;
        reg [4:0]               axi_w_cs, axi_w_ns;
        reg [LEN_W-1:0]         w_data_counter;
        reg [LEN_W-1:0]         user_w_len_ff;
        reg [ADDR_W-1:0]        user_w_addr_ff;
        reg [ASIZE_W-1:0]       user_w_awsize_ff;
        reg [ID_W-1:0]          user_w_awid_ff;
        reg                     ready_w_flag;
        reg                     start_w_ff;
        logic                    next_w_feed_in;
        logic                   burst_w_split_flag_ff;
        logic                   misalign_w_addr_flag_ff;
        logic [ADDR_W-1:0]      addr_w_tmp_ff;
        logic [LEN_W-1:0]       len_w_tmp_ff;
        logic [ADDR_W-1:0]      addr_w_split_tmp_ff;
        logic [LEN_W-1:0]       len_w_split_tmp_ff;
        logic [ADDR_W-1:0]      bytes_until_boundary;
        //logic [LEN_W-1:0]       beats_until_boundary;
        logic [ADDR_W-1:0]       beats_until_boundary;
        logic [LEN_W-1:0]       awlen_until_boundary;
        logic [3:0]             error_wrap;
        logic                   error_redux_or;
        logic                    no_beats_fit_flag;
        logic                    page_boundary_cross_no_split_flag;
        logic                    insufficient_wdata_flag;
        logic                    start_w_addr_misalign_flag;
        logic [3:0]             user_w_cmd_error_ff;
        logic                   underrun_flag_ff;

        logic [DATA_W-1:0]       w_data_final;
        logic [STRB_W-1:0]       w_strb_final;

        logic [LEN_W + DATA_W_BYTES_CLOG:0] total_bytes;
        logic [DATA_W_BYTES_CLOG-1:0] misalign_bytes;
        logic [LEN_W:0] beats_required;
        logic [LEN_W:0] len_decided;
        
        
// ---- FSM ---- //
        localparam WRITE_IDLE       = 'b00001;
        localparam WRITE_CHK_CMD    = 'b00010;
        localparam WRITE_ADDRESS    = 'b00100;
        localparam WRITE            = 'b01000;
        localparam WRITE_RESPONSE   = 'b10000;
    
        always_ff @ (posedge aclk)
        begin
            if(~aresetn)
            begin
                axi_w_cs <= WRITE_IDLE;
            end
        
            else
            begin
                axi_w_cs <= axi_w_ns;
            end
        end

        always_comb
        begin
            case(axi_w_cs)
            WRITE_IDLE:
            begin
                if(start_write)  axi_w_ns = WRITE_CHK_CMD;
                else             axi_w_ns = WRITE_IDLE;
            end

            WRITE_CHK_CMD:
            begin
                if(~error_redux_or) axi_w_ns = WRITE_ADDRESS;
                else                axi_w_ns = WRITE_IDLE;
            end
            
            WRITE_ADDRESS:
            begin
                if(m_axi_awready)   axi_w_ns = WRITE;
                else                axi_w_ns = WRITE_ADDRESS;
            end
        
            WRITE:
            begin
                if((w_data_counter == len_w_tmp_ff) && m_axi_wready)
                begin
                    axi_w_ns = WRITE_RESPONSE;
                end
            
                else
                begin
                    axi_w_ns = WRITE;
                end
            end
        
            WRITE_RESPONSE:
            begin
                if(m_axi_bvalid)
                begin
                    if(start_write) axi_w_ns = WRITE_CHK_CMD;
                    else            axi_w_ns = WRITE_IDLE;
                end
                else axi_w_ns = WRITE_RESPONSE;
            end
        
            default: axi_w_ns = WRITE_IDLE;
            endcase
        end

        assign next_w_feed_in       = (((axi_w_cs == WRITE_RESPONSE) && (m_axi_bvalid)) || (axi_w_cs == WRITE_IDLE)) ? 1 : 0;
        assign user_w_free          = (((axi_w_ns == WRITE_RESPONSE) || (axi_w_ns == WRITE_IDLE)) && ~start_w_ff && ~burst_w_split_flag_ff) ? 1 : 0;

        always_comb
        begin
            m_axi_awvalid  = 'h0;
            m_axi_awlen    = 'h0;
            m_axi_awlock   = 'h0;
            m_axi_awqos    = 'h0;
            m_axi_awregion = 'h0;
            m_axi_awaddr   = 'h0;
            m_axi_awprot   = 'h0;
            m_axi_awsize   = 'h0;
            m_axi_awburst  = 'b10;
            m_axi_awcache  = 'h0;
            m_axi_awid     = 'h0;
            m_axi_wvalid   = 'h0;
            m_axi_wdata    = 'h0;
            m_axi_wstrb    = 'h0;
            m_axi_wlast    = 'h0;
            m_axi_bready   = 'h0;
            //user_w_data_pop_req = 'h0;
            user_w_wready = 'h0;
            user_w_bid = 'h0;
            user_w_status = 'h0;
            user_w_bvalid = 'h0;

            if(axi_w_cs==WRITE_ADDRESS)
            begin
                m_axi_awvalid = 'h1;
                m_axi_awlen   = len_w_tmp_ff;
                m_axi_awaddr  = addr_w_tmp_ff;
                m_axi_awsize  = user_w_awsize_ff;
                m_axi_awid    = user_w_awid_ff;
            end

            w_data_final = (MISALIGN_ADJUST==0) ? user_w_data : aligned_w_data_final;
            w_strb_final = (MISALIGN_ADJUST==0) ? user_w_strb : aligned_w_strb_final;

            if(axi_w_cs==WRITE)
            begin
                case(BURST_POLICY)
                    0: 
                    begin
                        m_axi_wvalid  = 1; // data was pre-checked so no need to stall
                        m_axi_wdata   = w_data_final;
                        m_axi_wstrb   = w_strb_final;
                    end
                    
                    1: 
                    begin
                        //m_axi_wvalid  = ~(user_w_data_fifo_empty); // stall and wait if fifo is empty
                        m_axi_wvalid  = user_w_wvalid;
                        m_axi_wdata   = w_data_final;
                        m_axi_wstrb   = w_strb_final;
                    end

                    2: 
                    begin
                        m_axi_wvalid  = 1; // never stall, if fifo is empty then output dummy data
                        m_axi_wdata   = (~(user_w_data_fifo_empty)) ? w_data_final : 'h0;
                        m_axi_wstrb   = (~(user_w_data_fifo_empty)) ? w_strb_final : 'h0;
                    end
                endcase

                m_axi_wlast   = (w_data_counter == len_w_tmp_ff);
                //user_w_data_pop_req = (m_axi_wready && m_axi_wvalid && ~(user_w_data_fifo_empty));
                user_w_wready = m_axi_wready;
            end

            if(axi_w_cs == WRITE_RESPONSE)
            begin
                //m_axi_bready  = 'h1;
                m_axi_bready  = user_w_bready; // from fifo (ack)
                user_w_bvalid = m_axi_bvalid; // to fifo (req)

                user_w_bid    = m_axi_bid;
                user_w_status = m_axi_bresp;
            end
        end

// ---- Misaligned Address ---- //
    // TODO
    reg  [DATA_W_BYTES_CLOG-1:0]    w_addr_offset_ff;

    //reg carry_valid_ff;
    reg [DATA_W-1:0] carry_w_data_ff;
    reg [STRB_W-1:0] carry_w_strb_ff;

    logic [DATA_W-1:0] aligned_w_data;
    logic [DATA_W-1:0] carry_w_data;
    logic [DATA_W-1:0] aligned_w_data_final;
    logic [STRB_W-1:0] aligned_w_strb;
    logic [STRB_W-1:0] carry_w_strb;
    logic [STRB_W-1:0] aligned_w_strb_final;

    logic [DATA_W_CLOG-1:0] w_data_shift_left;
    logic [DATA_W_CLOG-1:0] w_data_shift_right;

    logic [STRB_W_CLOG-1:0] w_strb_shift_left;
    logic [STRB_W_CLOG-1:0] w_strb_shift_right;

    // Requirement:
        // - sequential logic for holding carry out data
            // carry valid (check wstrb bits)
            // carry data AND strb (flop the right-shifted signals for use in the next beat)
        // - combinational logic for w_data input shifting
            // shift data AND strb left (this becomes the data to use)
            // shift data AND strb right (this becomes the carry out)

            // aligned data + strb out that goes to the axi signals

    // EX:
        // 1. find the address offset + increase len -> len + 1
            // - detect if split burst is required (cross page boundary and/or len+1 > MAX_BURST_LEN)
        // 2. use the address offset to calculate:
            // - carry_out = (write data >> (address offset*8))
            // - data_to_use = (write data << (address offset*8))
        // 3. flop the carry out + write "data_to_use" to the w_data axi signal
            // flop : carry_out_ff <= carry_out
            // comb : m_axi_wdata = carry_out_ff | data_to_use;
        // 4. wlast
            // -> if split burst then we are required to carry data + wstrb  over to the next burst
            // -> if not:
                // comb : m_axi_wdata = carry_out_ff | 'h0;

        always_comb
        begin
            w_data_shift_left = (w_addr_offset_ff * BYTE);
            w_data_shift_right = (DATA_W - w_data_shift_left);

            w_strb_shift_left = (w_addr_offset_ff);
            w_strb_shift_right = (DATA_W_BYTES - w_strb_shift_left);

            if(w_addr_offset_ff == 0)
            begin
                aligned_w_data  =  user_w_data;
                carry_w_data    =  'h0;
                aligned_w_strb  =  user_w_strb;
                carry_w_strb    =  'h0;
            end

            else
            begin
                aligned_w_data  =  (user_w_data << (w_data_shift_left));
                carry_w_data    =  (user_w_data >> (w_data_shift_right));

                aligned_w_strb  =  (user_w_strb << (w_strb_shift_left));
                carry_w_strb    =  (user_w_strb >> (w_strb_shift_right));
            end
        end

// aligner
        logic                  align_carry_valid_ff;
        logic [DATA_W-1:0]     align_carry_w_data_ff;
        logic [DATA_W/8-1:0]   align_carry_w_strb_ff;

        always_ff @(posedge aclk) 
        begin
        if (~aresetn) 
        begin
            align_carry_valid_ff <= 1'b0;
            align_carry_w_data_ff <= '0;
            align_carry_w_strb_ff <= '0;
        end

        else if (start_w_ff && burst_w_split_flag_ff) 
        begin
            align_carry_valid_ff <= split_carry_valid_ff;  // burst start after split
            align_carry_w_data_ff <= split_carry_w_data_ff;
            align_carry_w_strb_ff <= split_carry_w_strb_ff;
        end

        else if (start_w_ff && ~burst_w_split_flag_ff) 
        begin
            align_carry_valid_ff <= 1'b0;  // reset at burst start
            align_carry_w_data_ff <= '0;
            align_carry_w_strb_ff <= '0;
        end

        else if (axi_w_cs==WRITE && m_axi_wready && m_axi_wvalid) 
        begin
            align_carry_valid_ff <= (|carry_w_strb);  // your shifted_lo leftover
            align_carry_w_data_ff <= carry_w_data;    // low bits that didn't fit
            align_carry_w_strb_ff <= carry_w_strb;
        end
    end

// splitter
        logic                  split_carry_valid_ff;
        logic [DATA_W-1:0]     split_carry_w_data_ff;
        logic [DATA_W/8-1:0]   split_carry_w_strb_ff;

        always_ff @(posedge aclk) 
        begin
            if (~aresetn) 
            begin
                split_carry_valid_ff <= 1'b0;
                split_carry_w_data_ff <= '0;
                split_carry_w_strb_ff <= '0;
            end

            else if ((axi_w_cs == WRITE) && m_axi_wvalid && m_axi_wready && m_axi_wlast && burst_w_split_flag_ff) 
            begin
                split_carry_valid_ff <= |carry_w_strb;
                split_carry_w_data_ff <= carry_w_data;
                split_carry_w_strb_ff <= carry_w_strb;
            end

            else if (start_w_ff && ~burst_w_split_flag_ff) 
            begin
                split_carry_valid_ff <= 'h0;  // burst start after split
                split_carry_w_data_ff <= 'h0;
                split_carry_w_strb_ff <= 'h0;
            end
        end

        always_comb
        begin
            aligned_w_data_final = 'h0;
            aligned_w_strb_final = 'h0;

            aligned_w_data_final = ((align_carry_valid_ff) ? align_carry_w_data_ff : 'h0)| aligned_w_data;
            aligned_w_strb_final = ((align_carry_valid_ff) ? align_carry_w_strb_ff : 'h0)| aligned_w_strb;

            // need to save the 'carry_w_data_ff' and 'carry_w_strb_ff' if 'burst_w_split_flag_ff' flag is set
        end

// ---- Underrun flag ---- //
        always_ff @ (posedge aclk)
        begin
            if(~aresetn)
            begin
                underrun_flag_ff <= 'h0;
            end

            else
            begin
                case(BURST_POLICY)
                0:
                begin
                    underrun_flag_ff <= 'h0;
                end

                1,2:
                begin
                    if(start_w_ff)
                    begin
                        underrun_flag_ff <= 'h0;
                    end

                    else if((axi_w_cs==WRITE) && (user_w_data_fifo_empty) && m_axi_wready && m_axi_wvalid)
                    begin
                        underrun_flag_ff <= 'h1;
                    end
                end
                endcase
            end
        end

        assign user_w_underrun_event = underrun_flag_ff;

// ---- Start + 1-stage pipeline + automatic start for cmd boundary split mechanism ---- //
        assign start_write  = (~error_redux_or) & start_w_ff;

        always_ff @ (posedge aclk)
        begin
            if(~aresetn)
            begin
                ready_w_flag          <= 1;
                start_w_ff            <= 0;

                user_w_len_ff           <= 0;
                user_w_addr_ff          <= 0;
                user_w_awsize_ff        <= 0;
                user_w_awid_ff          <= 0;

                w_addr_offset_ff        <= 'h0;
            end
            
            else
            begin
                if(ready_w_flag)
                begin
                    // TODO: misaligned address causes a split burst (1. across boundary, 2. len+1 > MAX_BURST_LEN, 3. both)

                    if((SPLIT_PAGE_BOUNDARY > 0) && burst_w_split_flag_ff)
                    begin
                        ready_w_flag      <= 0;
                        start_w_ff        <= 1;

                    end

                    else if(user_w_start)
                    begin
                        ready_w_flag      <= 0;
                        start_w_ff        <= 1;

                        user_w_len_ff     <= user_w_len;
                        user_w_addr_ff    <= user_w_addr;
                        user_w_awsize_ff  <= user_w_awsize;
                        user_w_awid_ff    <= user_w_awid;

                        w_addr_offset_ff  <= user_w_addr[DATA_W_BYTES_CLOG-1:0];
                    end
                end
                
                else if(next_w_feed_in & start_w_ff)
                begin
                    ready_w_flag      <= 1;
                    start_w_ff        <= 0;
                end
            end
        end
        
//---- Burst write beat counter for FSM ----//
        always_ff @ (posedge aclk)
        begin
            if(axi_w_cs == WRITE_IDLE || axi_w_cs == WRITE_RESPONSE) w_data_counter <= 'h0;
            
            else if(axi_w_cs == WRITE && m_axi_wready && m_axi_wvalid)//w_data_counter < len_w_tmp_ff)
            begin
                w_data_counter <= w_data_counter + 1'b1;
            end
            
            else w_data_counter <= w_data_counter;
        end

//---- Write status flop ----//
/*
        reg [RESP_W-1:0] user_w_status_ff;
        reg [ID_W-1:0]   user_w_bid_ff;

        assign user_w_status = user_w_status_ff;
        assign user_w_bid = user_w_bid_ff;

        always_ff (posedge aclk)
        begin
            if(~aresetn)
            begin
                user_w_status_ff  <= 'h0;
                user_w_bid_ff     <= 'h0;
            end

            else 
            begin
                if(start_w_ff)
                begin
                    user_w_status_ff  <= 'h0;
                    user_w_bid_ff     <= 'h0;
                end

                if(m_axi_bready && m_axi_bvalid)
                begin
                    user_w_status_ff  <= m_axi_bresp;
                    user_w_bid_ff     <= m_axi_bid;
                end
            end
        end
*/

//---- COMB + SEQ logic used for basis of error-checking and splitting bursts ----//
        always_comb
        begin
        // misaligned address
            total_bytes = ((user_w_len_ff + 1) << DATA_W_BYTES_CLOG);
            misalign_bytes = user_w_addr_ff[DATA_W_BYTES_CLOG-1:0];
            beats_required = ((total_bytes + misalign_bytes) + (DATA_W_BYTES-1)) >> DATA_W_BYTES_CLOG;

        // burst splitting
            // bytes until boundary
            bytes_until_boundary = PAGE_SIZE_BYTES - (user_w_addr_ff[PAGE_SIZE_BYTES_CLOG-1:0]);
            // burst beats until boundary
            beats_until_boundary = ((bytes_until_boundary + misalign_bytes) >> DATA_W_BYTES_CLOG);
            // adjusted for awlen (len-1)
            awlen_until_boundary = (beats_until_boundary == 0) ? 0 : beats_until_boundary-1;

        // error detection
            no_beats_fit_flag                   = (beats_until_boundary == 0);
            page_boundary_cross_no_split_flag   = (awlen_until_boundary < (beats_required-1));
            insufficient_wdata_flag             = (user_w_data_fifo_cnt < beats_required);
            start_w_addr_misalign_flag          = (misalign_bytes != 0);

            error_wrap = {
                            (MISALIGN_ADJUST == 0) && start_w_addr_misalign_flag, 
                            (BURST_POLICY == 0) && insufficient_wdata_flag, 
                            (SPLIT_PAGE_BOUNDARY == 0) && page_boundary_cross_no_split_flag,
                            no_beats_fit_flag
                        };

            error_redux_or = |error_wrap;

        // len decision
            len_decided = (page_boundary_cross_no_split_flag) ? awlen_until_boundary : ((beats_required > (MAX_BURST_BEATS-1)) ? MAX_BURST_BEATS-1 : user_w_len_ff);
            
        end

        always_ff @ (posedge aclk)
        begin
            if(~aresetn)
            begin
                addr_w_tmp_ff   <= 'h0;
                len_w_tmp_ff    <= 'h0;

                addr_w_split_tmp_ff     <= 'h0;
                len_w_split_tmp_ff      <= 'h0;
                burst_w_split_flag_ff   <= 'h0;

                misalign_w_addr_flag_ff <= 'h0;
            end

            else
            begin
                if(next_w_feed_in)
                begin
                    if(~burst_w_split_flag_ff)
                    begin

                        addr_w_tmp_ff   <= user_w_addr_ff & ~(DATA_W_BYTES-1);
                        len_w_tmp_ff    <= len_decided - 1;

                        if(SPLIT_PAGE_BOUNDARY > 0)
                        begin
                            if(beats_required > len_decided)
                            begin
                                burst_w_split_flag_ff     <= 1'b1;
                                addr_w_split_tmp_ff       <= user_w_addr_ff + (len_decided * DATA_W_BYTES) - misalign_bytes;
                                len_w_split_tmp_ff        <= (beats_required - len_decided) - 1;
                            end

                            else
                            begin
                                burst_w_split_flag_ff   <= 1'b0;
                                addr_w_split_tmp_ff     <= 'h0;
                                len_w_split_tmp_ff      <= 'h0;
                            end
                        end
                    end

                    else
                    begin
                        addr_w_tmp_ff   <= addr_w_split_tmp_ff;
                        len_w_tmp_ff    <= len_w_split_tmp_ff;

                        if(start_w_ff)
                        begin
                            burst_w_split_flag_ff   <= 1'b0;
                        end
                    end
                end
            end
        end

// ---- Error Flop set and clr for output port ----//
        assign user_w_cmd_error     = user_w_cmd_error_ff;

        always_ff @ (posedge aclk)
        begin
            if(~aresetn)
            begin
                user_w_cmd_error_ff <= 'h0;
            end

            else
            begin
                if(start_w_ff)
                begin
                    user_w_cmd_error_ff <= 'h0;
                end

                else if(axi_w_cs==WRITE_CHK_CMD)
                begin
                    user_w_cmd_error_ff <= error_wrap;
                end
            end
        end
    end
endgenerate

// AXI R ---------------------------------------------------
generate
    if(READ_EN)
    begin
        // FSM
        localparam READ_IDLE       = 5'b00001;
        localparam READ_ADDRESS    = 5'b00010;
        localparam READ_RESPONSE   = 5'b00100;

        logic start_read;
        
        reg [5:0] axi_r_cs, axi_r_ns;
    
        always @ (posedge aclk)
        begin
            if(~aresetn)
            begin
                axi_r_cs <= READ_IDLE;
            end
        
            else
            begin
                axi_r_cs <= axi_r_ns;
            end
        end

        always @ (*)
        begin
            case(axi_r_cs)
            READ_IDLE:
            begin
                if(start_read)  axi_r_ns = READ_ADDRESS;
                else            axi_r_ns = READ_IDLE;
            end
            
            READ_ADDRESS:
            begin
                if(m_axi_arready)  axi_r_ns = READ_RESPONSE;
                else               axi_r_ns = READ_ADDRESS;
            end

            READ_RESPONSE:
            begin
                if(m_axi_rlast)
                begin
                    if(start_read)  axi_r_ns = READ_ADDRESS;
                    else            axi_r_ns = READ_IDLE;
                end
            
                else
                begin
                    axi_r_ns = READ_RESPONSE;
                end
            end
        
            default: axi_r_ns = READ_IDLE;
            endcase
        end

        // System for locking-in next operation via flops
        reg [8-1:0]                 user_r_len_ff;
        reg [ADDR_W-1:0]            user_r_addr_ff;
        
        reg                         ready_r_flag;
        reg                         start_r_ff;
        logic                        next_r_feed_in;

        assign start_read = start_r_ff;

        always @ (posedge aclk)
        begin
            if(~aresetn)
            begin
                ready_r_flag            <= 1;
                start_r_ff              <= 0;
                //
                user_r_len_ff           <= 0;
                user_r_addr_ff          <= 0;
            end
            
            else
            begin
                if(ready_r_flag & user_r_start)
                begin
                    ready_r_flag      <= 0;
                    start_r_ff        <= 1;
                    //
                    user_r_len_ff     <= user_r_len;
                    user_r_addr_ff    <= user_r_addr;
                end
                
                else if(next_r_feed_in & start_r_ff)
                begin
                    ready_r_flag      <= 1;
                    start_r_ff        <= 0;
                end
            end
        end
        
        assign next_r_feed_in        = (((axi_r_cs == READ_RESPONSE) && (m_axi_rlast)) || (axi_r_cs == READ_IDLE)) ? 1 : 0;
        assign user_r_free           = (((axi_r_ns == READ_RESPONSE) || (axi_r_ns == READ_IDLE)) && ~start_r_ff) ? 1 : 0;
        // System for locking-in next operation via flops ^^^

        // AXI IN/OUT Signals
        /*
        always @ (posedge aclk)
        begin
            if(~aresetn)
            begin
                user_r_status_ff   <= 0;
            end
            
            else if(m_axi_rready && m_axi_rvalid)
            begin
                user_r_status_ff   <= m_axi_rresp;
            end

            else
            begin
                user_r_status_ff   <= 0;
            end
        end

        assign user_r_status         = user_r_status_ff;
        */
        
        assign user_r_status = 0;

        always_comb
        begin
            m_axi_arvalid   = 'h0;
            m_axi_arlen     = 'h0;
            m_axi_araddr    = 'h0;
            m_axi_rready    = 'h0;
            user_r_data     = 'h0;
            user_r_data_push_req = 'h0;

            if(axi_r_cs==READ_ADDRESS)
            begin
                m_axi_araddr      = user_r_addr_ff;
                m_axi_arlen       = user_r_len_ff;
                m_axi_arvalid     = 'h1;
            end
            
            if(axi_r_cs==READ_RESPONSE)
            begin
                m_axi_rready            = ~(user_r_fifo_full);
                user_r_data             = m_axi_rdata;
                user_r_data_push_req    = m_axi_rvalid && m_axi_rready;
            end
        end
    end
    
    else
    begin
        always_comb
        begin
            m_axi_araddr = 'h0;    // read address
            m_axi_arprot = 'h0;    // protection - privilege and securit level of transaction
            m_axi_arvalid = 'h0;   // 
            m_axi_arsize = 'h0;    //3'b100, // burst beat size - size of each transfer in the burst 3'b100 for 16 bytes/ 128 bit
            m_axi_arburst = 'h0;   // fixed burst = 00, incremental = 01, wrapped burst = 10
            m_axi_arcache = 'h0;   // cache type - how transaction interacts with caches
            m_axi_arlen = 'h0;     // number of data transfers in the burst (0-255) (done)
            m_axi_arlock = 'h0;    // lock type - indicates if transaction is part of locked sequence
            m_axi_arqos = 'h0;     // quality of service - transaction indication of priority level
            m_axi_arregion = 'h0;  // region identifier - identifies targetted region
            m_axi_arid = 'h0;
            m_axi_rready = 'h0;    // read ready - 0 = not ready, 1 = ready
        end
    end
endgenerate
endmodule
